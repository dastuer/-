library verilog;
use verilog.vl_types.all;
entity div_fre_test is
end div_fre_test;
