library verilog;
use verilog.vl_types.all;
entity BDPSK_test is
end BDPSK_test;
