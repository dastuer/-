library verilog;
use verilog.vl_types.all;
entity dif_encoder_test is
end dif_encoder_test;
