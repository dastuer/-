library verilog;
use verilog.vl_types.all;
entity PN_Seq_test is
end PN_Seq_test;
